`ifndef _AXI_REG_FILE_DEF_H_
`define _AXI_REG_FILE_DEF_H_

// `include "axi_reg_file.svh"
// 
// `define MEMORY_MAPPED       1'b1
// `define NO_MEMORY_MAPPED    1'b0
// `define TRIGGER_ON_WRITE    1'b1
// `define NO_TRIGGER_ON_WRITE 1'b0
// `define CLEAR_ON_READ       1'b1
// `define NO_CLEAR_ON_READ    1'b0
// 
// typedef struct packed {
//     logic   [`AXI_REG_FILE_ADDR_WIDTH-1:0]  addr;
//     logic   [31:0]                          val;
//     logic                                   memory_mapped;
//     logic                                   trigger_on_write;
//     logic                                   clear_on_read;
// } reg_entry_t;

`endif
